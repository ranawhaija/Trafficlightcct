CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
770 80 1364 707
42991634 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 308 555 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
6666 0 0
2
5.89624e-315 0
0
13 Logic Switch~
5 247 552 0 1 11
0 16
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9365 0 0
2
5.89624e-315 0
0
13 Logic Switch~
5 491 31 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3251 0 0
2
5.89624e-315 0
0
13 Logic Switch~
5 442 37 0 1 11
0 21
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5481 0 0
2
5.89624e-315 0
0
13 Logic Switch~
5 32 118 0 1 11
0 23
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7788 0 0
2
5.89624e-315 0
0
13 Logic Switch~
5 85 94 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3273 0 0
2
5.89624e-315 0
0
13 Logic Switch~
5 132 84 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3761 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 231 194 0 1 2
10 3
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 919 424 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4244 0 0
2
5.89624e-315 0
0
9 2-In NOR~
219 856 393 0 3 22
0 5 6 4
0
0 0 624 270
6 74LS02
-21 -24 21 -16
3 U8B
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5225 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 917 355 0 1 2
10 6
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
768 0 0
2
5.89624e-315 0
0
5 7415~
219 791 358 0 4 22
0 9 8 7 6
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 5 0
1 U
5735 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 917 296 0 1 2
10 5
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5881 0 0
2
5.89624e-315 0
0
5 7415~
219 792 299 0 4 22
0 9 8 10 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
3275 0 0
2
5.89624e-315 0
0
9 2-In NOR~
219 836 199 0 3 22
0 12 13 11
0
0 0 624 270
6 74LS02
-21 -24 21 -16
3 U8A
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4203 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 916 230 0 1 2
10 11
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 915 166 0 1 2
10 13
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9102 0 0
2
5.89624e-315 0
0
14 Logic Display~
6 917 102 0 1 2
10 12
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5586 0 0
2
5.89624e-315 0
0
5 7415~
219 780 170 0 4 22
0 9 10 14 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
525 0 0
2
5.89624e-315 0
0
5 7415~
219 779 108 0 4 22
0 15 14 7 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
6206 0 0
2
5.89624e-315 0
0
5 7474~
219 599 365 0 6 22
0 17 18 3 17 10 7
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 1 0
1 U
3418 0 0
2
5.89624e-315 0
0
6 74LS74
17 603 191 0 12 25
0 3 20 17 17 3 19 17 17 15
9 8 14
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 0 1 0 0 0
1 U
9312 0 0
2
5.89624e-315 0
0
7 74LS153
119 397 346 0 14 29
0 26 10 10 10 15 8 27 28 29
30 21 21 18 31
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
7419 0 0
2
5.89624e-315 0
0
7 74LS153
119 398 192 0 14 29
0 32 10 7 16 15 8 33 16 10
7 21 21 20 19
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
472 0 0
2
5.89624e-315 0
0
7 Pulser~
4 37 294 0 10 12
0 34 35 22 36 0 0 5 5 3
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4714 0 0
2
5.89624e-315 0
0
7 74LS190
134 181 207 0 14 29
0 24 22 2 23 23 23 23 23 3
37 38 39 40 41
0
0 0 4848 0
7 74LS190
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9386 0 0
2
5.89624e-315 0
0
61
3 1 2 0 0 8320 0 26 6 0 0 3
143 198
85 198
85 106
1 0 3 0 0 8320 0 8 0 0 4 3
215 198
215 110
364 110
1 9 3 0 0 128 0 8 26 0 0 2
215 198
219 198
0 1 3 0 0 4096 0 0 22 0 0 4
356 110
522 110
522 155
571 155
1 3 4 0 0 8320 0 9 10 0 0 3
903 428
903 426
862 426
1 0 5 0 0 4096 0 10 0 0 12 2
871 374
871 300
2 0 6 0 0 4096 0 10 0 0 8 2
853 374
853 359
4 1 6 0 0 8320 0 12 11 0 0 3
812 358
812 359
901 359
0 3 7 0 0 8192 0 0 12 24 0 3
681 329
681 367
767 367
0 2 8 0 0 4096 0 0 12 14 0 3
728 299
728 358
767 358
0 1 9 0 0 4096 0 0 12 15 0 3
739 290
739 349
767 349
4 1 5 0 0 8320 0 14 13 0 0 3
813 299
813 300
901 300
0 3 10 0 0 8192 0 0 14 21 0 3
756 309
756 308
768 308
0 2 8 0 0 12288 0 0 14 37 0 4
656 277
707 277
707 299
768 299
0 1 9 0 0 4224 0 0 14 23 0 3
718 173
718 290
768 290
3 1 11 0 0 8320 0 15 16 0 0 3
842 232
842 234
900 234
1 0 12 0 0 4096 0 15 0 0 20 2
851 180
851 108
2 0 13 0 0 4096 0 15 0 0 19 2
833 180
833 170
1 4 13 0 0 4224 0 17 19 0 0 2
899 170
801 170
1 4 12 0 0 8320 0 18 20 0 0 3
901 106
901 108
800 108
2 0 10 0 0 4096 0 19 0 0 33 3
756 170
756 364
629 364
3 0 14 0 0 4096 0 19 0 0 25 2
756 179
679 179
10 1 9 0 0 0 0 22 19 0 0 4
641 173
743 173
743 161
756 161
0 3 7 0 0 8192 0 0 20 34 0 4
656 329
692 329
692 117
755 117
12 2 14 0 0 8320 0 22 20 0 0 4
641 218
679 218
679 108
755 108
1 0 15 0 0 4096 0 20 0 0 39 2
755 99
656 99
2 0 10 0 0 0 0 23 0 0 33 2
365 319
282 319
3 0 10 0 0 0 0 23 0 0 33 2
365 328
282 328
4 0 10 0 0 0 0 23 0 0 33 2
365 337
282 337
8 0 16 0 0 4096 0 24 0 0 35 2
366 219
248 219
9 0 10 0 0 0 0 24 0 0 33 2
366 228
282 228
10 0 7 0 0 0 0 24 0 0 34 2
366 237
298 237
5 2 10 0 0 8320 0 21 24 0 0 5
629 347
629 416
282 416
282 165
366 165
6 3 7 0 0 12416 0 21 24 0 0 6
623 329
656 329
656 430
298 430
298 174
366 174
4 1 16 0 0 8320 0 24 2 0 0 3
366 183
248 183
248 539
0 6 8 0 0 4096 0 0 24 37 0 3
347 277
347 201
366 201
11 6 8 0 0 12416 0 22 23 0 0 6
635 209
656 209
656 277
347 277
347 355
365 355
0 5 15 0 0 4096 0 0 23 39 0 3
329 192
329 346
365 346
9 5 15 0 0 12416 0 22 24 0 0 6
635 164
656 164
656 58
329 58
329 192
366 192
5 0 3 0 0 0 0 22 0 0 41 2
571 200
517 200
0 3 3 0 0 4224 0 0 21 4 0 3
517 153
517 347
575 347
0 4 17 0 0 4224 0 0 21 44 0 3
549 227
549 377
599 377
7 1 17 0 0 0 0 22 21 0 0 3
565 218
565 302
599 302
0 8 17 0 0 0 0 0 22 46 0 3
549 182
549 227
565 227
3 7 17 0 0 0 0 22 22 0 0 2
565 173
565 218
0 4 17 0 0 0 0 0 22 47 0 3
549 43
549 182
565 182
3 1 17 0 0 0 0 22 3 0 0 3
565 173
565 43
491 43
13 2 18 0 0 8320 0 23 21 0 0 3
429 328
429 329
575 329
14 6 19 0 0 4224 0 24 22 0 0 4
430 219
545 219
545 209
571 209
13 2 20 0 0 4224 0 24 22 0 0 4
430 174
504 174
504 164
571 164
0 12 21 0 0 4096 0 0 23 52 0 3
442 310
442 391
435 391
0 11 21 0 0 0 0 0 23 53 0 3
442 237
442 310
435 310
0 12 21 0 0 4096 0 0 24 54 0 3
442 155
442 237
436 237
1 11 21 0 0 4224 0 4 24 0 0 3
442 49
442 156
436 156
2 3 22 0 0 8320 0 26 25 0 0 4
149 189
105 189
105 285
61 285
0 8 23 0 0 8320 0 0 26 57 0 3
32 234
32 243
149 243
0 7 23 0 0 0 0 0 26 58 0 3
32 225
32 234
149 234
0 6 23 0 0 0 0 0 26 59 0 3
32 216
32 225
149 225
5 0 23 0 0 0 0 26 0 0 60 3
149 216
32 216
32 207
1 4 23 0 0 0 0 5 26 0 0 3
32 130
32 207
149 207
1 1 24 0 0 4224 0 7 26 0 0 3
132 96
132 180
143 180
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
934 88 971 112
944 96 960 112
2 G1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
929 154 966 178
939 162 955 178
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
933 215 970 239
943 223 959 239
2 R1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
930 283 967 307
940 291 956 307
2 G2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
935 342 972 366
945 350 961 366
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
940 407 977 431
950 415 966 431
2 R2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
